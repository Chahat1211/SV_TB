interface inf;
	logic[1:0] a;
	logic[1:0] b;
 	logic[1:0] c;
	logic[1:0] d;
	logic[1:0] sel;
	logic[1:0] out;
endinterface
	
