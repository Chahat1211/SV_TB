interface inf (input logic clk);
	logic d;
	logic reset;
	logic q;
endinterface
